// Language: VHDL
// Type: Unit Converter
// Category: Hardware
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
