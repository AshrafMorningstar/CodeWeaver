// Language: VHDL
// Type: CLI Calculator
// Category: Hardware
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
