// Language: VHDL
// Type: Simple Encryption/Decryption
// Category: Hardware
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
