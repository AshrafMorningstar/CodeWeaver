// Language: VHDL
// Type: Number Guessing Game
// Category: Hardware
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
