// Language: VHDL
// Type: File Processor
// Category: Hardware
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
print('Line {i}');
